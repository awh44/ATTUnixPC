library ieee;
use ieee.std_logic_1164.all;

package types is
	type bus_array is array(natural range <>) of std_logic_vector(0 downto 0);
end types;
